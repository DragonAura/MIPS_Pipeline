`timescale 1ns / 1ns

module testCPU(

    );

    reg clk, rst;
    // wire [31:0] memAddr;
    // wire [31:0] deviceData;
    // wire [31:0] memOut;
    reg rx;
    wire tx;
    wire [6:0] leds;
    wire [3:0] ano;
    wire dot;
    // wire led;

    wire memRead, memWrite;

    wire [31:0] memAddr;
    wire [31:0] memData;
    wire [31:0] deviceData;


    CPU cpu(
            .clk(clk),
            .rst(rst),
            .memRead_MEM(memRead),
            .memWrite_MEM(memWrite),
            .memAddr(memAddr),
            .memDat(memData),
            .deviceData(deviceData)
        );

    LED led(
            .clk(clk),
            .rst(rst),
            .memWrite(memWrite),
            .dataIn(memData),
            .address(memAddr),
            .digi({ano, dot, leds})
        );

    UART uart(
             .clk(clk),
             .rst(rst),
             .rx(rx),
             .memRead(memRead),
             .memWrite(memWrite),
             .dataIn(memData),
             .address(memAddr),
             .uartData(deviceData),
             .tx(tx)
         );

    // top topmodule(clk, rst, rx, tx, leds, ano, dot);


    integer i, j;
    wire [31:0] data0, data1, data2, data3, data4, data5, data6, data7, data8, data9, data10, num;
    assign data0 = 32'h00000000;
    assign data1 = 32'h00000001;
    assign data2 = 32'h00000002;
    assign data3 = 32'h00000003;
    assign data4 = 32'h00000004;
    assign data5 = 32'h00000005;
    assign data6 = 32'h00000006;
    assign data7 = 32'h00000007;
    assign data8 = 32'h00000008;
    assign data9 = 32'h00000009;
    assign data10 = 32'hffffffff;
    assign num = 20;

    initial begin
        clk = 0;
        rst = 0;
        rx = 1;
        #2 rst = 1;
        #2 rst = 0;
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = num[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data10[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data7[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data6[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data1[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data3[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data4[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data5[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data8[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data9[8 * i + j];
            end
            #100 rx = 1;
        end
        for (i = 3; i >= 0; i = i - 1) begin
            #100 rx = 0;
            for (j = 0; j < 8; j = j + 1) begin
                #100 rx = data0[8 * i + j];
            end
            #100 rx = 1;
        end

    end

    always #5 clk = ~clk;

endmodule
